interface basic_if
    integer a;
    integer b;
endinterface