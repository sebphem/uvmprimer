import uvm_pkg::*;

class quarter_uvm_agent extends uvm_agent;
    //register with the factory
    `uvm_component_utils(quarter_uvm_agent);

    //add in the 
    uvm_analysis_port#()
endclass