import uvm_pkg::*;
module tb;
    




endmodule