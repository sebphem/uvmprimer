import uvm_pkg::*;


interface quarter_if;
    logic clk;
    logic reset_n;
    logic quarter_slot;
    logic ticket;
endinterface

