class basic_cov

    


endclass