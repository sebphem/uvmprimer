module scoreboard(
    bfm
);
    
endmodule