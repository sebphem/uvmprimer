import uvm_pkg::*;

class basic_test extends uvm_test;

    `uvm_component_utils(basic_test);
    basic_env env;

    function new(string name="basic_test",uvm_component parent)

endclass